LIBRARY ieee;
USE ieee. std_logic_1164.all;
 
ENTITY relogio_digital IS
	PORT(CLEAR: IN BIT;
	     CLOCK: IN STD_LOGIC;
	  MIN, SEG: OUT BIT_VECTOR(3 DOWNTO 0));
END relogio_digital;

 
ARCHITECTURE arch OF relogio_digital IS

COMPONENT cont_mod10 IS
	PORT(CLEAR: IN BIT;
		 CLOCK: IN STD_LOGIC;
	       SEG: OUT BIT_VECTOR(3 DOWNTO 0));
END COMPONENT;

SIGNAL Q, QM: BIT_VECTOR(3 DOWNTO 0) := "0000";
SIGNAL QB, QBM: BIT_VECTOR(3 DOWNTO 0) := "1111";

BEGIN
	contador_segundos: cont_mod10 PORT MAP(CLEAR, CLOCK, SEG);

	--FFM0: JK_FF PORT MAP(QBM(1) OR QBM(2), '1'           , CLEAR, CLOCK, QM(0), QBM(0));
	--FFM1: JK_FF PORT MAP(QBM(0) AND QM(2), QM(0) OR QM(2), CLEAR, CLOCK, QM(1), QBM(1));
	--FFM2: JK_FF PORT MAP(QM(0)  AND QM(1), QM(0) OR QM(1), CLEAR, CLOCK, QM(2), QBM(2));
END arch;
