LIBRARY ieee;
USE ieee. std_logic_1164.all;
 
ENTITY cont_mod6 IS
	PORT(CLEAR: IN BIT;
		 CLOCK: IN STD_LOGIC;
	    OUTPUT: OUT BIT_VECTOR(3 DOWNTO 0));
END cont_mod6;

 
ARCHITECTURE arch OF cont_mod6 IS

COMPONENT JK_FF IS
	PORT(J,K,CLEAR: IN BIT;
	         CLOCK: IN STD_LOGIC;
	         Q, QB: OUT BIT);
END COMPONENT;

SIGNAL Q: BIT_VECTOR(3 DOWNTO 0) := "0000";
SIGNAL QB: BIT_VECTOR(3 DOWNTO 0) := "1111";

BEGIN
	FFM0: JK_FF PORT MAP(QB(1) OR QB(2), '1'         , CLEAR, CLOCK, Q(0), QB(0));
	FFM1: JK_FF PORT MAP(Q(0) AND QB(2), Q(0) OR Q(2), CLEAR, CLOCK, Q(1), QB(1));
	FFM2: JK_FF PORT MAP(Q(0)  AND Q(1), Q(0) OR Q(1), CLEAR, CLOCK, Q(2), QB(2));
	
	OUTPUT(0) <= Q(0);
	OUTPUT(1) <= Q(1);
	OUTPUT(2) <= Q(2);
	OUTPUT(3) <= Q(3);
END arch;